
module SSDNiosSoftwareEmbarcado (
	clk_clk,
	medidordesempenho_conduit_readdata,
	reset_reset_n);	

	input		clk_clk;
	output	[31:0]	medidordesempenho_conduit_readdata;
	input		reset_reset_n;
endmodule
